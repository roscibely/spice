*Base comum tjb
v1 1 0 dc 5V
R1 1 2 1000
Q1 2 0 3 npnt
.model npnt npn(Is=1.8104e-15 Bf=50)
v2 3 0 dc 1V
.control 
dc v1 0 5V 1V
dc v2 0 1V 1V
plot v(2)
.endc
.END 
